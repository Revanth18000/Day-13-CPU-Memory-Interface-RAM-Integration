module simple_ram (
    input clk,
    input we,
    input [3:0] addr,
    input [7:0] data_in,
    output reg [7:0] data_out
);

    reg [7:0] mem [0:15];

    always @(posedge clk) begin
        if (we)
            mem[addr] <= data_in;     // WRITE
        else
            data_out <= mem[addr];   // READ
    end

endmodule